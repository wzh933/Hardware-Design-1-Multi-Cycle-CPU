`timescale 1ps / 1ps
`include "alu.v"
module st3_exe (  // ִ��
    input EXE_valid,  // ִ�м���Ч�ź�
    input [149:0] ID_EXE_bus_r,  //ID->EXE����
    output EXE_over,
    output [105:0] EXE_MEM_bus,  //EXE->MEM����

    // չʾpc
    output [31:0] EXE_pc
);
  // ID->EXE���� begin
  // EXE��Ҫ�õ�����Ϣ
  // ALU����Դ�������Ϳ����ź�
  wire [11:0] alu_control;
  wire [31:0] alu_operand1;
  wire [31:0] alu_operand2;

  // �´���Ҫ�õ��� load / store ��Ϣ
  wire [3:0] mem_control;  // MEM��Ҫʹ�õĿ����ź�
  wire [31:0] store_data;  // store�����Ĵ������

  // д����Ҫ�õ�����Ϣ
  wire rf_wen;
  wire [4:0] rf_wdest;

  // pc
  wire [31:0] pc;
  assign  {alu_control, alu_operand1, alu_operand2, mem_control, store_data, rf_wen, rf_wdest, pc} = ID_EXE_bus_r;
  //ID->EXE end

  // ALU begin
  wire [31:0] alu_result;

  // ����aluģ��
  alu alu_module (
      .alu_control(alu_control),  // input, 12, ALU�����ź�
      .alu_src1(alu_operand1),  // input, 32, ALU������1
      .alu_src2(alu_operand2),  // input, 32, ALU������2
      .alu_result(alu_result)  // output, 32, ALU���
  );
  // ALU end

  // EXEִ����� begin
  // �����Ƕ����ڵģ��������������
  // ������ALU���㶼����һ�������
  // ��EXEģ��һ�ľ���������в���
  // ��EXE_valid����EXE_over�ź�
  assign EXE_over = EXE_valid;
  // EXEִ����� end

  // EXE->MEM���� begin
  assign EXE_MEM_bus = {
    mem_control,
    store_data,  // load / store ��Ϣ��store����
    alu_result,  // ALU������ 
    rf_wen,
    rf_wdest,  // WB��Ҫʹ�õ��ź�
    pc  // pcֵ
  };
  // EXE->MEM���� end

  // display EXE_pc begin
  assign EXE_pc = pc;
  // display EXE_pc end
endmodule
